/****************************************************************************************
*****************************************************************************************
Name: 
	PCEn
	
Description: 
	

Subject:
	Microprocessors Design - ITESO

Author:
	Cesar Carlos Robles Martinez 

Date:
	14/04/2019
*****************************************************************************************
*****************************************************************************************/

module PCEn

//Input ports 
(
	input Branch,
	input PCWrite,

//Output ports 

	output PCEn_out
);

/*******************************************************************************
*												CODE  															
*******************************************************************************/

assign PCEn_out = Branch | PCWrite; 

endmodule
